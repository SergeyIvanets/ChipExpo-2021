`timescale 1ns/1ps
// add latency
`define PIPELINE 

// no latency
//`define NOPIPELINE
